-- megafunction wizard: %ALTLVDS%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altlvds_tx 

-- ============================================================
-- File Name: alt_lvds_tx.vhd
-- Megafunction Name(s):
-- 			altlvds_tx
--
-- Simulation Library Files(s):
-- 			altera_mf
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 8.0 Build 215 05/29/2008 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2008 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY altera_mf;
USE altera_mf.all;

ENTITY alt_lvds_tx IS
	PORT
	(
		tx_in		: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
		tx_inclock		: IN STD_LOGIC  := '0';
		tx_out		: OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
		tx_outclock		: OUT STD_LOGIC 
	);
END alt_lvds_tx;


ARCHITECTURE SYN OF alt_lvds_tx IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire1	: STD_LOGIC ;



	COMPONENT altlvds_tx
	GENERIC (
		common_rx_tx_pll		: STRING;
		deserialization_factor		: NATURAL;
		implement_in_les		: STRING;
		inclock_data_alignment		: STRING;
		inclock_period		: NATURAL;
		inclock_phase_shift		: NATURAL;
		intended_device_family		: STRING;
		lpm_type		: STRING;
		number_of_channels		: NATURAL;
		outclock_alignment		: STRING;
		outclock_divide_by		: NATURAL;
		outclock_phase_shift		: NATURAL;
		outclock_resource		: STRING;
		output_data_rate		: NATURAL;
		registered_input		: STRING;
		use_external_pll		: STRING
	);
	PORT (
			tx_out	: OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
			tx_outclock	: OUT STD_LOGIC ;
			tx_in	: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
			tx_inclock	: IN STD_LOGIC 
	);
	END COMPONENT;

BEGIN
	tx_out    <= sub_wire0(1 DOWNTO 0);
	tx_outclock    <= sub_wire1;

	altlvds_tx_component : altlvds_tx
	GENERIC MAP (
		common_rx_tx_pll => "OFF",
		deserialization_factor => 8,
		implement_in_les => "OFF",
		inclock_data_alignment => "UNUSED",
		inclock_period => 8000,
		inclock_phase_shift => 0,
		intended_device_family => "Stratix II",
		lpm_type => "altlvds_tx",
		number_of_channels => 2,
		outclock_alignment => "UNUSED",
		outclock_divide_by => 1,
		outclock_phase_shift => 0,
		outclock_resource => "AUTO",
		output_data_rate => 750,
		registered_input => "TX_CORECLK",
		use_external_pll => "OFF"
	)
	PORT MAP (
		tx_in => tx_in,
		tx_inclock => tx_inclock,
		tx_out => sub_wire0,
		tx_outclock => sub_wire1
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: Clock_Choices STRING "TX_CORECLK"
-- Retrieval info: PRIVATE: Clock_Mode NUMERIC "0"
-- Retrieval info: PRIVATE: Data_rate STRING "750"
-- Retrieval info: PRIVATE: Deser_Factor NUMERIC "8"
-- Retrieval info: PRIVATE: Enable_DPA_Mode STRING "OFF"
-- Retrieval info: PRIVATE: Ext_PLL STRING "OFF"
-- Retrieval info: PRIVATE: INCLOCK_PHASE_SHIFT STRING "0.00"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Stratix II"
-- Retrieval info: PRIVATE: Int_Device STRING "Stratix II"
-- Retrieval info: PRIVATE: LVDS_Mode NUMERIC "0"
-- Retrieval info: PRIVATE: Le_Serdes STRING "OFF"
-- Retrieval info: PRIVATE: Num_Channel NUMERIC "2"
-- Retrieval info: PRIVATE: OUTCLOCK_PHASE_SHIFT STRING "0.00"
-- Retrieval info: PRIVATE: Outclock_Divide_By NUMERIC "1"
-- Retrieval info: PRIVATE: PLL_Enable NUMERIC "0"
-- Retrieval info: PRIVATE: PLL_Freq STRING "125.00"
-- Retrieval info: PRIVATE: PLL_Period STRING "8.000"
-- Retrieval info: PRIVATE: Reg_InOut NUMERIC "1"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: PRIVATE: Use_Clock_Resc STRING "AUTO"
-- Retrieval info: PRIVATE: Use_Common_Rx_Tx_Plls NUMERIC "0"
-- Retrieval info: PRIVATE: Use_CoreClock NUMERIC "0"
-- Retrieval info: PRIVATE: Use_Lock NUMERIC "0"
-- Retrieval info: PRIVATE: Use_Pll_Areset NUMERIC "0"
-- Retrieval info: PRIVATE: Use_Tx_Out_Phase NUMERIC "1"
-- Retrieval info: CONSTANT: COMMON_RX_TX_PLL STRING "OFF"
-- Retrieval info: CONSTANT: DESERIALIZATION_FACTOR NUMERIC "8"
-- Retrieval info: CONSTANT: IMPLEMENT_IN_LES STRING "OFF"
-- Retrieval info: CONSTANT: INCLOCK_DATA_ALIGNMENT STRING "UNUSED"
-- Retrieval info: CONSTANT: INCLOCK_PERIOD NUMERIC "8000"
-- Retrieval info: CONSTANT: INCLOCK_PHASE_SHIFT NUMERIC "0"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Stratix II"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "altlvds_tx"
-- Retrieval info: CONSTANT: NUMBER_OF_CHANNELS NUMERIC "2"
-- Retrieval info: CONSTANT: OUTCLOCK_ALIGNMENT STRING "UNUSED"
-- Retrieval info: CONSTANT: OUTCLOCK_DIVIDE_BY NUMERIC "1"
-- Retrieval info: CONSTANT: OUTCLOCK_PHASE_SHIFT NUMERIC "0"
-- Retrieval info: CONSTANT: OUTCLOCK_RESOURCE STRING "AUTO"
-- Retrieval info: CONSTANT: OUTPUT_DATA_RATE NUMERIC "750"
-- Retrieval info: CONSTANT: REGISTERED_INPUT STRING "TX_CORECLK"
-- Retrieval info: CONSTANT: USE_EXTERNAL_PLL STRING "OFF"
-- Retrieval info: USED_PORT: tx_in 0 0 16 0 INPUT NODEFVAL tx_in[15..0]
-- Retrieval info: USED_PORT: tx_inclock 0 0 0 0 INPUT_CLK_EXT GND tx_inclock
-- Retrieval info: USED_PORT: tx_out 0 0 2 0 OUTPUT NODEFVAL tx_out[1..0]
-- Retrieval info: USED_PORT: tx_outclock 0 0 0 0 OUTPUT NODEFVAL tx_outclock
-- Retrieval info: CONNECT: @tx_in 0 0 16 0 tx_in 0 0 16 0
-- Retrieval info: CONNECT: tx_out 0 0 2 0 @tx_out 0 0 2 0
-- Retrieval info: CONNECT: @tx_inclock 0 0 0 0 tx_inclock 0 0 0 0
-- Retrieval info: CONNECT: tx_outclock 0 0 0 0 @tx_outclock 0 0 0 0
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: GEN_FILE: TYPE_NORMAL alt_lvds_tx.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL alt_lvds_tx.ppf TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL alt_lvds_tx.inc TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL alt_lvds_tx.cmp FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL alt_lvds_tx.bsf TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL alt_lvds_tx_inst.vhd FALSE
-- Retrieval info: LIB_FILE: altera_mf
