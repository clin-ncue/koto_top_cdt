module GenTrigger(clk,rst,ene,ntrig,gap,trigger);

input wire clk;
input wire rst;
input wire ene;
input wire [15:0] ntrig;
input wire [7:0] gap;

output reg trigger;

//reg [7:0] gap_reg;
reg [7:0] counter;
reg [15:0] ntrig_reg;

always @( posedge clk)
begin

//	gap_reg = gap - 1'b1;

	if
	(rst)
	begin
		ntrig_reg = 16'b0;
		counter = 8'b0;
	end

	if( ene && ntrig_reg <= ntrig )
	begin
		if(counter==gap)
		begin
			trigger = 1'b1;
			ntrig_reg = ntrig_reg + 1'b1;
			counter = 8'b0;
		end
		else 
		begin
			trigger = 1'b0;
		end
		counter = counter + 1'b1;
	end
	else
	begin
		trigger = 1'b0;
	end

	
end

endmodule