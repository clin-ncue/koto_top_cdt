-- megafunction wizard: %ALTLVDS%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altlvds_tx 

-- ============================================================
-- File Name: CL_ALTLVDS_Tx_1.vhd
-- Megafunction Name(s):
-- 			altlvds_tx
--
-- Simulation Library Files(s):
-- 			altera_mf
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 9.1 Build 350 03/24/2010 SP 2 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2010 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY altera_mf;
USE altera_mf.all;

ENTITY CL_ALTLVDS_Tx_1 IS
	PORT
	(
		pll_areset		: IN STD_LOGIC  := '0';
		tx_in		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		tx_inclock		: IN STD_LOGIC  := '0';
		tx_out		: OUT STD_LOGIC_VECTOR (0 DOWNTO 0)
	);
END CL_ALTLVDS_Tx_1;


ARCHITECTURE SYN OF cl_altlvds_tx_1 IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (0 DOWNTO 0);



	COMPONENT altlvds_tx
	GENERIC (
		common_rx_tx_pll		: STRING;
		deserialization_factor		: NATURAL;
		implement_in_les		: STRING;
		inclock_data_alignment		: STRING;
		inclock_period		: NATURAL;
		inclock_phase_shift		: NATURAL;
		intended_device_family		: STRING;
		lpm_hint		: STRING;
		lpm_type		: STRING;
		number_of_channels		: NATURAL;
		outclock_resource		: STRING;
		output_data_rate		: NATURAL;
		registered_input		: STRING;
		use_external_pll		: STRING
	);
	PORT (
			pll_areset	: IN STD_LOGIC ;
			tx_out	: OUT STD_LOGIC_VECTOR (0 DOWNTO 0);
			tx_in	: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
			tx_inclock	: IN STD_LOGIC 
	);
	END COMPONENT;

BEGIN
	tx_out    <= sub_wire0(0 DOWNTO 0);

	altlvds_tx_component : altlvds_tx
	GENERIC MAP (
		common_rx_tx_pll => "ON",
		deserialization_factor => 8,
		implement_in_les => "OFF",
		inclock_data_alignment => "UNUSED",
		inclock_period => 32000,
		inclock_phase_shift => 1000,
		intended_device_family => "Stratix II",
		lpm_hint => "CBX_MODULE_PREFIX=CL_ALTLVDS_Tx_1",
		lpm_type => "altlvds_tx",
		number_of_channels => 1,
		outclock_resource => "AUTO",
		output_data_rate => 250,
		registered_input => "TX_CLKIN",
		use_external_pll => "OFF"
	)
	PORT MAP (
		pll_areset => pll_areset,
		tx_in => tx_in,
		tx_inclock => tx_inclock,
		tx_out => sub_wire0
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: Clock_Choices STRING "TX_CLKIN"
-- Retrieval info: PRIVATE: Clock_Mode NUMERIC "1"
-- Retrieval info: PRIVATE: Data_rate STRING "250"
-- Retrieval info: PRIVATE: Deser_Factor NUMERIC "8"
-- Retrieval info: PRIVATE: Enable_DPA_Mode STRING "OFF"
-- Retrieval info: PRIVATE: Ext_PLL STRING "OFF"
-- Retrieval info: PRIVATE: INCLOCK_PHASE_SHIFT STRING "90.00"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Stratix II"
-- Retrieval info: PRIVATE: Int_Device STRING "Stratix II"
-- Retrieval info: PRIVATE: LVDS_Mode NUMERIC "0"
-- Retrieval info: PRIVATE: Le_Serdes STRING "OFF"
-- Retrieval info: PRIVATE: Num_Channel NUMERIC "1"
-- Retrieval info: PRIVATE: OUTCLOCK_PHASE_SHIFT STRING "0"
-- Retrieval info: PRIVATE: Outclock_Divide_By NUMERIC "2"
-- Retrieval info: PRIVATE: PLL_Enable NUMERIC "0"
-- Retrieval info: PRIVATE: PLL_Freq STRING "31.25"
-- Retrieval info: PRIVATE: PLL_Period STRING "32.000"
-- Retrieval info: PRIVATE: Reg_InOut NUMERIC "1"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: PRIVATE: Use_Clock_Resc STRING "AUTO"
-- Retrieval info: PRIVATE: Use_Common_Rx_Tx_Plls NUMERIC "1"
-- Retrieval info: PRIVATE: Use_CoreClock NUMERIC "0"
-- Retrieval info: PRIVATE: Use_Lock NUMERIC "0"
-- Retrieval info: PRIVATE: Use_Pll_Areset NUMERIC "1"
-- Retrieval info: PRIVATE: Use_Tx_Out_Phase NUMERIC "1"
-- Retrieval info: CONSTANT: COMMON_RX_TX_PLL STRING "ON"
-- Retrieval info: CONSTANT: DESERIALIZATION_FACTOR NUMERIC "8"
-- Retrieval info: CONSTANT: IMPLEMENT_IN_LES STRING "OFF"
-- Retrieval info: CONSTANT: INCLOCK_DATA_ALIGNMENT STRING "UNUSED"
-- Retrieval info: CONSTANT: INCLOCK_PERIOD NUMERIC "32000"
-- Retrieval info: CONSTANT: INCLOCK_PHASE_SHIFT NUMERIC "1000"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Stratix II"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "altlvds_tx"
-- Retrieval info: CONSTANT: NUMBER_OF_CHANNELS NUMERIC "1"
-- Retrieval info: CONSTANT: OUTCLOCK_RESOURCE STRING "AUTO"
-- Retrieval info: CONSTANT: OUTPUT_DATA_RATE NUMERIC "250"
-- Retrieval info: CONSTANT: REGISTERED_INPUT STRING "TX_CLKIN"
-- Retrieval info: CONSTANT: USE_EXTERNAL_PLL STRING "OFF"
-- Retrieval info: USED_PORT: pll_areset 0 0 0 0 INPUT GND pll_areset
-- Retrieval info: USED_PORT: tx_in 0 0 8 0 INPUT NODEFVAL tx_in[7..0]
-- Retrieval info: USED_PORT: tx_inclock 0 0 0 0 INPUT_CLK_EXT GND tx_inclock
-- Retrieval info: USED_PORT: tx_out 0 0 1 0 OUTPUT NODEFVAL tx_out[0..0]
-- Retrieval info: CONNECT: @tx_in 0 0 8 0 tx_in 0 0 8 0
-- Retrieval info: CONNECT: tx_out 0 0 1 0 @tx_out 0 0 1 0
-- Retrieval info: CONNECT: @tx_inclock 0 0 0 0 tx_inclock 0 0 0 0
-- Retrieval info: CONNECT: @pll_areset 0 0 0 0 pll_areset 0 0 0 0
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: GEN_FILE: TYPE_NORMAL CL_ALTLVDS_Tx_1.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL CL_ALTLVDS_Tx_1.ppf TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL CL_ALTLVDS_Tx_1.inc TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL CL_ALTLVDS_Tx_1.cmp FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL CL_ALTLVDS_Tx_1.bsf TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL CL_ALTLVDS_Tx_1_inst.vhd FALSE
-- Retrieval info: LIB_FILE: altera_mf
-- Retrieval info: CBX_MODULE_PREFIX: ON
