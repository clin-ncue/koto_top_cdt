-- megafunction wizard: %PARALLEL_ADD%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: parallel_add 

-- ============================================================
-- File Name: CL_ADDER_4x1.vhd
-- Megafunction Name(s):
-- 			parallel_add
--
-- Simulation Library Files(s):
-- 			altera_mf
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 9.1 Build 350 03/24/2010 SP 2 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2010 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY altera_mf;
USE altera_mf.altera_mf_components.all;

ENTITY CL_ADDER_4x1 IS
	PORT
	(
		data0x		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		data1x		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		data2x		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		data3x		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (2 DOWNTO 0)
	);
END CL_ADDER_4x1;


ARCHITECTURE SYN OF cl_adder_4x1 IS

--	type ALTERA_MF_LOGIC_2D is array (NATURAL RANGE <>, NATURAL RANGE <>) of STD_LOGIC;

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (2 DOWNTO 0);
	SIGNAL sub_wire1	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire2	: ALTERA_MF_LOGIC_2D (3 DOWNTO 0, 0 DOWNTO 0);
	SIGNAL sub_wire3	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire4	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire5	: STD_LOGIC_VECTOR (0 DOWNTO 0);

BEGIN
	sub_wire5    <= data0x(0 DOWNTO 0);
	sub_wire4    <= data1x(0 DOWNTO 0);
	sub_wire3    <= data2x(0 DOWNTO 0);
	result    <= sub_wire0(2 DOWNTO 0);
	sub_wire1    <= data3x(0 DOWNTO 0);
	sub_wire2(3, 0)    <= sub_wire1(0);
	sub_wire2(2, 0)    <= sub_wire3(0);
	sub_wire2(1, 0)    <= sub_wire4(0);
	sub_wire2(0, 0)    <= sub_wire5(0);

	parallel_add_component : parallel_add
	GENERIC MAP (
		msw_subtract => "NO",
		pipeline => 0,
		representation => "UNSIGNED",
		result_alignment => "LSB",
		shift => 0,
		size => 4,
		width => 1,
		widthr => 3,
		lpm_type => "parallel_add"
	)
	PORT MAP (
		data => sub_wire2,
		result => sub_wire0
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Stratix II"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: CONSTANT: MSW_SUBTRACT STRING "NO"
-- Retrieval info: CONSTANT: PIPELINE NUMERIC "0"
-- Retrieval info: CONSTANT: REPRESENTATION STRING "UNSIGNED"
-- Retrieval info: CONSTANT: RESULT_ALIGNMENT STRING "LSB"
-- Retrieval info: CONSTANT: SHIFT NUMERIC "0"
-- Retrieval info: CONSTANT: SIZE NUMERIC "4"
-- Retrieval info: CONSTANT: WIDTH NUMERIC "1"
-- Retrieval info: CONSTANT: WIDTHR NUMERIC "3"
-- Retrieval info: USED_PORT: data0x 0 0 1 0 INPUT NODEFVAL "data0x[0..0]"
-- Retrieval info: USED_PORT: data1x 0 0 1 0 INPUT NODEFVAL "data1x[0..0]"
-- Retrieval info: USED_PORT: data2x 0 0 1 0 INPUT NODEFVAL "data2x[0..0]"
-- Retrieval info: USED_PORT: data3x 0 0 1 0 INPUT NODEFVAL "data3x[0..0]"
-- Retrieval info: USED_PORT: result 0 0 3 0 OUTPUT NODEFVAL "result[2..0]"
-- Retrieval info: CONNECT: @data 1 3 1 0 data3x 0 0 1 0
-- Retrieval info: CONNECT: @data 1 2 1 0 data2x 0 0 1 0
-- Retrieval info: CONNECT: @data 1 1 1 0 data1x 0 0 1 0
-- Retrieval info: CONNECT: @data 1 0 1 0 data0x 0 0 1 0
-- Retrieval info: CONNECT: result 0 0 3 0 @result 0 0 3 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL CL_ADDER_4x1.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL CL_ADDER_4x1.inc TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL CL_ADDER_4x1.cmp FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL CL_ADDER_4x1.bsf TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL CL_ADDER_4x1_inst.vhd FALSE
-- Retrieval info: LIB_FILE: altera_mf
