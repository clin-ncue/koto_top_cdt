-- megafunction wizard: %Shift register (RAM-based)%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altshift_taps 

-- ============================================================
-- File Name: CL_Pipe_16x128.vhd
-- Megafunction Name(s):
-- 			altshift_taps
--
-- Simulation Library Files(s):
-- 			altera_mf
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 9.1 Build 350 03/24/2010 SP 2 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2010 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY altera_mf;
USE altera_mf.all;

ENTITY CL_Pipe_16x128 IS
	PORT
	(
		clock		: IN STD_LOGIC ;
		shiftin		: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
		shiftout		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		taps		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
	);
END CL_Pipe_16x128;


ARCHITECTURE SYN OF cl_pipe_16x128 IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (15 DOWNTO 0);
	SIGNAL sub_wire1	: STD_LOGIC_VECTOR (15 DOWNTO 0);



	COMPONENT altshift_taps
	GENERIC (
		lpm_hint		: STRING;
		lpm_type		: STRING;
		number_of_taps		: NATURAL;
		tap_distance		: NATURAL;
		width		: NATURAL
	);
	PORT (
			taps	: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
			clock	: IN STD_LOGIC ;
			shiftout	: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
			shiftin	: IN STD_LOGIC_VECTOR (15 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	taps    <= sub_wire0(15 DOWNTO 0);
	shiftout    <= sub_wire1(15 DOWNTO 0);

	altshift_taps_component : altshift_taps
	GENERIC MAP (
		lpm_hint => "RAM_BLOCK_TYPE=M512",
		lpm_type => "altshift_taps",
		number_of_taps => 1,
		tap_distance => 128,
		width => 16
	)
	PORT MAP (
		clock => clock,
		shiftin => shiftin,
		taps => sub_wire0,
		shiftout => sub_wire1
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: ACLR NUMERIC "0"
-- Retrieval info: PRIVATE: CLKEN NUMERIC "0"
-- Retrieval info: PRIVATE: GROUP_TAPS NUMERIC "0"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Stratix II"
-- Retrieval info: PRIVATE: NUMBER_OF_TAPS NUMERIC "1"
-- Retrieval info: PRIVATE: RAM_BLOCK_TYPE NUMERIC "0"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: PRIVATE: TAP_DISTANCE NUMERIC "128"
-- Retrieval info: PRIVATE: WIDTH NUMERIC "16"
-- Retrieval info: CONSTANT: LPM_HINT STRING "RAM_BLOCK_TYPE=M512"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "altshift_taps"
-- Retrieval info: CONSTANT: NUMBER_OF_TAPS NUMERIC "1"
-- Retrieval info: CONSTANT: TAP_DISTANCE NUMERIC "128"
-- Retrieval info: CONSTANT: WIDTH NUMERIC "16"
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL clock
-- Retrieval info: USED_PORT: shiftin 0 0 16 0 INPUT NODEFVAL shiftin[15..0]
-- Retrieval info: USED_PORT: shiftout 0 0 16 0 OUTPUT NODEFVAL shiftout[15..0]
-- Retrieval info: USED_PORT: taps 0 0 16 0 OUTPUT NODEFVAL taps[15..0]
-- Retrieval info: CONNECT: @shiftin 0 0 16 0 shiftin 0 0 16 0
-- Retrieval info: CONNECT: shiftout 0 0 16 0 @shiftout 0 0 16 0
-- Retrieval info: CONNECT: taps 0 0 16 0 @taps 0 0 16 0
-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: GEN_FILE: TYPE_NORMAL CL_Pipe_16x128.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL CL_Pipe_16x128.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL CL_Pipe_16x128.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL CL_Pipe_16x128.bsf TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL CL_Pipe_16x128_inst.vhd FALSE
-- Retrieval info: LIB_FILE: altera_mf
